
`timescale 1ns / 1ps
`default_nettype none

module main	(
  input wire CLOCK_50,            //On Board 50 MHz
  input wire [9:0] SW,            // On board Switches
  input wire [3:0] KEY,           // On board push buttons
  output wire [6:0] HEX0,         // HEX displays
  output wire [6:0] HEX1,
  output wire [6:0] HEX2,
  output wire [6:0] HEX3,
  output wire [6:0] HEX4,
  output wire [6:0] HEX5,
  output wire [9:0] LEDR,         // LEDs
  output wire [7:0] x,            // VGA pixel coordinates
  output wire [6:0] y,
  output wire [2:0] colour,       // VGA pixel colour (0-7)
  output wire plot,               // Pixel drawn when this is pulsed
  output wire vga_resetn          // VGA resets to black when this is pulsed (NOT CURRENTLY AVAILABLE)
);

  mux m1(LEDR,SW);

endmodule


module mux(LEDR, SW);
    input [9:0] SW;
    output [9:0] LEDR;

    mux2to1 u0(
        .x(SW[0]),
        .y(SW[1]),
        .s(SW[9]),
        .m(LEDR[0])
        );
endmodule

module mux2to1(x, y, s, m);
    input x; //select 0
    input y; //select 1
    input s; //select signal
    output m; //output

    //assign m = s & y | ~s & x;
    // OR
    assign m = s ? y : x;

endmodule
